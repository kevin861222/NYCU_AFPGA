module Lab8_0811127(input a , output b);

endmodule
